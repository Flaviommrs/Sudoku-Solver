LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE Sudoku  IS
	TYPE states_UC IS (FETCH, DECODE, EX);
	
	
	component bank IS
	GENERIC (
		WORDSIZE : NATURAL := 4
	);
	PORT (
		WR_EN, RD_EN,
		clear,
		clock		: IN 	STD_LOGIC;
		WR_ADDR,
		RD_ADDR1	: IN	STD_LOGIC_VECTOR (6 DOWNTO 0);
		DATA_IN		: IN	STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0);
		Player_in	: in std_logic;
		DATA_OUT1	: OUT	STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0);
		Player_out	: out std_logic;
	);
	END component;
	
	
	
	component BitmapVerifier is
	port(vecline, vecoluwn, vecregion: in std_logic_vector(8 downto 0);
		enable	: in std_logic;
		pos_x, pos_y: in std_logic_vector(3 downto 0);
		result:	out std_logic);
	end component;
	
	component bmap is
	port(
	pos_x, pos_y: in std_logic_vector(3 downto 0);
	clk, enable, clear: std_logic;
	x, y, region :out  std_logic_vector(8 downto 0)
  );
	end component;
	
	component count_adder IS
	GENERIC(modulo: Integer := 8);
	PORT(Clock: IN STD_LOGIC ;
	     E, Set, LOAD, CLEAR, signpositive: IN STD_LOGIC ;
         BCD: BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0) := (others =>'0');
         PAR_IN: in STD_LOGIC_VECTOR(3 DOWNTO 0);
         CARRY_OUT: out STD_LOGIC);
	END component ;
	
	component reg is
	GENERIC ( N : INTEGER ) ;
	port(data_in: in std_logic_vector(N-1 downto 0);
		 load, clear, clk: in std_logic;
		 player_in: in std_logic;
		 data_out: out std_logic_vector(N-1 downto 0);
		 player_out: in std_logic )
	end component;
	
	component Mux9to1 is
	port(vec1, vec2, vec3, vec4, vec5, vec6, vec7, vec8, vec9 : std_logic_vector(8 downto 0);
		 number: std_logic_vector(3 downto 0);
		 vec_out: std_logic_vector(8 downto 0)
		 );
	end component;
	
	component InputInterface is
	port(enter,
		 clear,
		 y,
	 	 x,
	 	 xdir,
	 	 ydir,
	 	 done: in std_logic;
	 	 data: in std_logic_vector(3 downto 0);
	 	 load,
	 	 go,
		 erase: out std_logic;
		 data_out: out std_logic_vector(3 downto 0);
	 	 positionX, positionY: out std_logic_vector(3 downto 0)
	 	);
	end component;
	
	
	
	
	
	
	
	
	
	
	
	
	
	COMPONENT memory IS
		GENERIC (
			WORDSIZE		: NATURAL	:= 8;
			BITS_OF_ADDR	: NATURAL	:= 16;
			MIF_FILE		: STRING	:= ""
		);
		PORT (
			clock   : IN	STD_LOGIC;
			we      : IN	STD_LOGIC;
			address : IN	STD_LOGIC_VECTOR(BITS_OF_ADDR-1 DOWNTO 0);
			datain  : IN	STD_LOGIC_VECTOR(WORDSIZE-1 DOWNTO 0);
			dataout : OUT	STD_LOGIC_VECTOR(WORDSIZE-1 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT reg IS
		GENERIC (
			WORDSIZE	: NATURAL := 32
		);
		PORT (
			clock,
			load,
			clear	: IN	STD_LOGIC;
			datain	: IN	STD_LOGIC_VECTOR(WORDSIZE-1 DOWNTO 0);
			dataout : OUT	STD_LOGIC_VECTOR(WORDSIZE-1 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT bank IS
		GENERIC (
			WORDSIZE : NATURAL := 32
		);
		PORT (
			WR_EN, RD_EN,
			clear,
			clock		: IN 	STD_LOGIC;
			WR_ADDR,
			RD_ADDR1,
			RD_ADDR2	: IN	STD_LOGIC_VECTOR (4 DOWNTO 0);
			DATA_IN		: IN	STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0);
			DATA_OUT1,
			DATA_OUT2	: OUT	STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT ALU IS
		GENERIC (
			WORDSIZE	: NATURAL := 4
		);
		PORT (
			A, B		: IN		STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0);
			Op			: IN		STD_LOGIC_VECTOR (1 DOWNTO 0);
			F			: BUFFER	STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0);
			Z, C, V, N	: OUT		STD_LOGIC
		);
	END COMPONENT;

	COMPONENT PC IS
		GENERIC (
			increment	: NATURAL := 4;
			WORDSIZE	: NATURAL := 32
		);
		PORT (
			clock,
			load,
			enable		: IN		STD_LOGIC;
			DATA_IN		: IN		STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0);
			DATA_OUT	: BUFFER	STD_LOGIC_VECTOR (WORDSIZE-1 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT UC IS
		PORT (
			clear,
			clock			: IN	STD_LOGIC;
			instruction		: IN	STD_LOGIC_VECTOR (2 DOWNTO 0);
			IR_Ld, PC_Inc, ALU_2_DBus, DM_Rd, DM_Wr, PC_Ld_En, Reg_2_IO, IO_2_Reg, Reg_Wr, Stat_Wr,
			DM_2_DBus		: OUT	STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT processor
		PORT (
			clock				:	 IN STD_LOGIC;
			reset				:	 IN STD_LOGIC;
			IO_IN				:	 IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			DBus				:	 OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			RSource1			:	 OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			RSource2			:	 OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			IO_OUT				:	 OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			IM_address			:	 OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			IM_instruction_out	:	 OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			instruction			:	 OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			stat_CVNZ			:	 OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Pc_Ld				:	 OUT STD_LOGIC;
			IR_Ld				:	 OUT STD_LOGIC;
			Pc_Inc				:	 OUT STD_LOGIC;
			ALU_2_DBus			:	 OUT STD_LOGIC;
			DM_Rd				:	 OUT STD_LOGIC;
			DM_Wr				:	 OUT STD_LOGIC;
			PC_Ld_En			:	 OUT STD_LOGIC;
			Reg_2_IO			:	 OUT STD_LOGIC;
			IO_2_Reg			:	 OUT STD_LOGIC;
			Reg_Wr				:	 OUT STD_LOGIC;
			Stat_Wr				:	 OUT STD_LOGIC;
			DM_2_DBus			:	 OUT STD_LOGIC
		);
	END COMPONENT;
	
	-- COMPONENTES ADICIONAIS PARA O nM
	component ram is
		generic(
			depth : natural := 12;
			width: natural := 32;
			init_file : string := ""
		);
		port(
			clk : in std_logic;
			memwrite:  in std_logic;
			ra, wa : in std_logic_vector(depth-1 downto 0);
			writedata : in std_logic_vector(width-1 downto 0);
			memdata : out std_logic_vector(width-1 downto 0)
		);
	end component;
	
	component rom is
		generic (
			depth : natural   := 32;
			width : natural   := 32; 
			init_file : string := ""
		);
		port(
		  clk : in std_logic;
		  adr: in std_logic_vector(depth-1 downto 0);
		  memdata: out std_logic_vector(width-1 downto 0)
	    );
	end component;
	
	component vga_text_mode is
		generic (
			init_file1 : string := "";
			init_file2 : string := ""
		);	
		port(
			clk : in std_logic;
			reset : in std_logic;
			write: in std_logic_vector(1 downto 0);
			showmem : in std_logic;
			wa : in std_logic_vector(11 downto 0);
			wd : in std_logic_vector(7 downto 0);
			HS : out std_logic;
			VS : out std_logic;
			blank : out std_logic;
			column : out std_logic_vector(6 downto 0);
			row : out std_logic_vector(5 downto 0);
			pixel : out std_logic
		);
	end component;
	
	component vga_timing is
		port(
			clk : in std_logic;
			reset : in std_logic;
			HS : out std_logic;
			VS : out std_logic;
			pixel_x : out std_logic_vector(9 downto 0);
			pixel_y : out std_logic_vector(9 downto 0);
			last_column : out std_logic;
			last_row : out std_logic;
			blank : out std_logic
		);
	end component;
	
	component flopar is
		generic(
			width: natural := 32
		);
		port(
			clk, reset: in std_logic;
			d: in  std_logic_vector(width-1 downto 0);
			q: out std_logic_vector(width-1 downto 0)
		);
	end component;
	
	component bin2hexascii is
		port(
			bin   : in std_logic_vector(3 downto 0);
			ascii : out std_logic_vector(7 downto 0)
		);
	end component;
	
	component m1ps2vga is
		port(
			clk : in std_logic;
			reset : in std_logic;
			start : in std_logic;
			pc, ir, dbus, rs1, rs2 : in std_logic_vector(31 downto 0); 
			stat : in std_logic_vector(3 downto 0);
			pcld, pcinc, irwr, regwr, statwr, dmwr, dmrd, dm2dbus,
				alu2dbus, reg2io, io2reg : in std_logic;
			aluop : in std_logic_vector(1 downto 0);
			memdata : in std_logic_vector(31 downto 0);
			regdata : in std_logic_vector(31 downto 0);
			
			vgawrite : out std_logic_vector(1 downto 0);
			vgawa : out std_logic_vector(11 downto 0);
			vgawd : out std_logic_vector(7 downto 0);
			memraddr : out std_logic_vector(7 downto 0);
			regaddr : out std_logic_vector(4 downto 0)
		);
	end component;
	
	component freqdiv is
		generic (DIV : natural := 2);
		port (
			clk : in std_logic;
			reset : in std_logic;
			clk_out : out std_logic
		);
	end component;
	
	component mM is
		generic(
			dm_init : string := ""
		);
		port(
			clk  : in std_logic;
			reset : in std_logic;
			pc, ir, dbus, rs1, rs2 : in std_logic_vector(31 downto 0);
			stat : in std_logic_vector(3 downto 0);
			pcld, pcinc, irwr, regwr, statwr, dmwr, dmrd, dm2dbus,
				alu2dbus, reg2io, io2reg : in std_logic;
			aluop : in std_logic_vector(1 downto 0);
			showscreen : in std_logic;
			vgaHS, vgaVS, vgablank, vgapixel : out std_logic;
			vgacolumn : out std_logic_vector(6 downto 0);
			vgarow : out std_logic_vector(5 downto 0)
			);
	end component;
	
	component counter is
		generic (
			nmax : natural := 128
		);
		port(	
			clk : in std_logic;
			reset : in std_logic;
			recount : in std_logic;
			encount : in std_logic;
			n : out natural range 0 to nmax;
			onmax : out std_logic
		);
	end component;
	
END PACKAGE;
